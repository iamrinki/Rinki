***** Spice Netlist for Cell 'lab9_inv' *****

************** Module lab9_inv **************
.subckt lab9_inv vin vout
m1 vout vin gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
m2 vout vin vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
.ends lab9_inv


