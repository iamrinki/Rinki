***** Spice Netlist for Cell 'lab10_inv' *****

************** Module lab10_inv **************
.subckt lab10_inv
m0 n0 n2 n1 n3 scmosn w='0.6u' l='0.4u' m='1' 
NULL scmosp4
NULL scmosp4
NULL scmosp4
.ends lab10_inv

************** Module scmosp4 **************
.subckt scmosp4
.ends scmosp4


.end

