magic
tech scmos
timestamp 1623394990
<< nwell >>
rect -26 1 34 22
<< ntransistor >>
rect 0 -13 2 -5
<< ptransistor >>
rect 0 8 2 16
<< ndiffusion >>
rect -5 -13 0 -5
rect 2 -13 13 -5
<< pdiffusion >>
rect -5 8 0 16
rect 2 8 13 16
<< ndcontact >>
rect -9 -13 -5 -5
rect 13 -13 17 -5
<< pdcontact >>
rect -9 8 -5 16
rect 13 8 17 16
<< psubstratepcontact >>
rect -19 -13 -15 -5
<< nsubstratencontact >>
rect -19 8 -15 16
<< polysilicon >>
rect 0 16 2 18
rect 0 5 2 8
rect 0 -5 2 1
rect 0 -15 2 -13
<< polycontact >>
rect -3 1 2 5
<< metal1 >>
rect -20 19 20 22
rect -15 8 -9 19
rect -5 2 -3 5
rect 13 -5 16 8
rect -15 -16 -9 -5
rect -20 -19 20 -16
<< labels >>
rlabel metal1 -15 21 -15 21 5 vdd!
rlabel metal1 -14 -18 -14 -18 1 gnd!
rlabel metal1 -5 4 -5 4 1 in!
rlabel metal1 13 4 13 4 1 out!
<< end >>
